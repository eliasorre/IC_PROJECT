* Pixel sensor
**********************************************************************
**        Copyright (c) 2021 Carsten Wulff Software, Norway
** *******************************************************************
** Created       : wulff at 2021-7-22
** *******************************************************************
**  The MIT License (MIT)
**
**  Permission is hereby granted, free of charge, to any person obtaining a copy
**  of this software and associated documentation files (the "Software"), to deal
**  in the Software without restriction, including without limitation the rights
**  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
**  copies of the Software, and to permit persons to whom the Software is
**  furnished to do so, subject to the following conditions:
**
**  The above copyright notice and this permission notice shall be included in all
**  copies or substantial portions of the Software.
**
**  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
**  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
**  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
**  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
**  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
**  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
**  SOFTWARE.
**
**********************************************************************

* Paramater
.param w_n = 0.09u
.param w_p = {w_n}
.param lu = 0.15u


.SUBCKT PIXEL_SENSOR VBN1 VRAMP VRESET ERASE EXPOSE READ
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS


XS1 VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR

XC1 VCMP_OUT VSTORE VRAMP VDD VSS VBN1 COMP

XM1 READ VCMP_OUT DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY

.ENDS

.SUBCKT MEMORY READ VCMP_OUT
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

XM1 VCMP_OUT DATA_0 READ VSS MEMCELL
XM2 VCMP_OUT DATA_1 READ VSS MEMCELL
XM3 VCMP_OUT DATA_2 READ VSS MEMCELL
XM4 VCMP_OUT DATA_3 READ VSS MEMCELL
XM5 VCMP_OUT DATA_4 READ VSS MEMCELL
XM6 VCMP_OUT DATA_5 READ VSS MEMCELL
XM7 VCMP_OUT DATA_6 READ VSS MEMCELL
XM8 VCMP_OUT DATA_7 READ VSS MEMCELL

.ENDS

.SUBCKT MEMCELL CMP DATA READ VSS
M1 VG CMP DATA VSS nmos  w=1u  l=0.13u
M2 DATA READ DMEM VSS nmos  w=0.2u  l=0.13u
M3 DMEM VG VSS VSS nmos  w=1u  l=0.13u
C1 VG VSS 1p
.ENDS

.SUBCKT SENSOR VRESET VSTORE ERASE EXPOSE VDD VSS

* * Capacitor to model gate-source capacitance
C1 VSTORE VSS 100f
Rleak VSTORE VSS 100T

* Switch to reset voltage on capacitor
MR VRESET ERASE VSTORE VSTORE nmos w=0.13u l=0.65u 
* Switch to expose pixel
ME VSTORE EXPOSE VPG VPG nmos w=0.13u l=0.65u 

* Model photocurrent
Rphoto VPG VSS 1G
.ENDS

.SUBCKT COMP VCMP_OUT VSTORE VRAMP VDD VSS VBN1

MP1 MPS1 MPS1 VDD VDD pmos w=w_p l=lu m=12
MP2 MPS2 MPS1 VDD VDD pmos w=w_p l=lu m=12

** The diff-pair of transistors, set to moderate inversion
MN3 MPS1 VSTORE MNS3 MNS3 nmos w=w_n l=lu
MN4 MPS2 VRAMP MNS3 MNS3 nmos w=w_n l=lu 

** Cascade Current Mirror to drive the diff-amp and gain-inverter
XCUR MNS3 MP6S VSS CASCADE_CURRENT_MIRROR

MP6 MP6S MPS2 VDD VDD pmos w=w_p l=lu m=12
*XCUR2 MP6S VSS CASCADE_CURRENT_MIRROR

** Inverter
MP8 VCMP_OUT MP6S VDD VDD pmos w=w_p l=lu m=12
MN9 VCMP_OUT MP6S VSS VSS nmos w=w_n l=lu m=5 

.ENDS

.SUBCKT CASCADE_CURRENT_MIRROR VIN1 VIN2 VOUT 
Isource VOUT MN2D dc 1u  
MN1 MN1D MN1D VOUT VOUT nmos w=(w_n*2.5) l=lu m=5
MN2 MN2D MN2D MN1D MN1D nmos w=(w_n*2.5) l=lu m=5

// Make two identical contact points, two drive two different parts of the circuit
MNO11 MNO12D MN1D VOUT VOUT nmos w=(w_n*2.5) l=lu m=25
MNO12 VIN1 MN2D MNO12D MNO12D nmos w=(w_n*2.5) l=lu m=25

MNO21 MNO22D MN1D VOUT VOUT nmos w=(w_n *2.5) l=lu m=25
MNO22 VIN2 MN2D MNO22D MNO22D nmos w=(w_n*2.5) l=lu m=25
.ENDS
