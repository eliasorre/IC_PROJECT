* Pixel sensor
**********************************************************************
**        Copyright (c) 2021 Carsten Wulff Software, Norway
** *******************************************************************
** Created       : wulff at 2021-7-22
** *******************************************************************
**  The MIT License (MIT)
**
**  Permission is hereby granted, free of charge, to any person obtaining a copy
**  of this software and associated documentation files (the "Software"), to deal
**  in the Software without restriction, including without limitation the rights
**  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
**  copies of the Software, and to permit persons to whom the Software is
**  furnished to do so, subject to the following conditions:
**
**  The above copyright notice and this permission notice shall be included in all
**  copies or substantial portions of the Software.
**
**  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
**  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
**  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
**  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
**  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
**  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
**  SOFTWARE.
**
**********************************************************************

* Paramater
.param w_n = 0.65
.param w_p = {w_n * 2.57}
.param lu = 0.13u


.SUBCKT PIXEL_SENSOR VBN1 VRAMP VRESET ERASE EXPOSE READ
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS


XS1 VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR

XC1 VCMP_OUT VSTORE VRAMP VDD VSS VBN1 COMP

XM1 READ VCMP_OUT DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY

.ENDS

.SUBCKT CASCADE_CURRENT_MIRROR VDD VSS 

Isource VSS MN3D dc 1u  

MN1 MN1D MN1D VSS VSS nmos w=w l=l m=5
MN2 MN2D MN1D VSS VSS nmos w=w l=l m=25
MN3 MN3D MN3D MN1D MN1D nmos w=w l=l m=5
MN4 VDD MN3D MN2D MN2D nmos w=w l=l m=25



.SUBCKT MEMORY READ VCMP_OUT
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

XM1 VCMP_OUT DATA_0 READ VSS MEMCELL
XM2 VCMP_OUT DATA_1 READ VSS MEMCELL
XM3 VCMP_OUT DATA_2 READ VSS MEMCELL
XM4 VCMP_OUT DATA_3 READ VSS MEMCELL
XM5 VCMP_OUT DATA_4 READ VSS MEMCELL
XM6 VCMP_OUT DATA_5 READ VSS MEMCELL
XM7 VCMP_OUT DATA_6 READ VSS MEMCELL
XM8 VCMP_OUT DATA_7 READ VSS MEMCELL

.ENDS

.SUBCKT MEMCELL CMP DATA READ VSS
M1 VG CMP DATA VSS nmos  w=0.2u  l=0.13u
M2 DATA READ DMEM VSS nmos  w=0.4u  l=0.13u
M3 DMEM VG VSS VSS nmos  w=1u  l=0.13u
C1 VG VSS 1p
.ENDS

.SUBCKT SENSOR VRESET VSTORE ERASE EXPOSE VDD VSS

MN9 MN9S VPG MN9S VSS nmos w=w_n l=lu
MN10 MN9S EXPOSE VSTORE VSS nmos w=w_n l=lu
MN11 VSS VSTORE VSS VSS nmos w=w_n l=lu
MN12 VRESET ERASE VSTORE VSS nmos w=w_n l=lu

* C1 VSTORE VSS 100f
* Rleak VSTORE VSS 100T   

* Model photocurrent
* Rphoto VPG VSS 1G
.ENDS

.SUBCKT COMP VCMP_OUT VSTORE VRAMP VDD VSS VBN1

MP1 VDD MPS1 MPS1 VSS pmos w=w_p l=lu
MP2 VDD MPS1 MPS2 VSS pmos w=w_p l=lu
MN3 MPS1 VSTORE MNS3 VSS nmos w=w_n l=lu
MN4 MPS2 VRAMP MNS3 VSS nmos w=w_n l=lu
MN5 MNS3 VBN1 VSS VSS nmos w=w_n l=lu
MP6 VDD MPS2 MP6S VSS pmos w=w_p l=lu
MN7 MP6S VBN1 VSS VSS nmos w=w_n l=lu
MP8 VDD MP6S VCMP_OUT VSS pmos w=w_p l=lu
MN9 VCMP_OUT MP6S VSS VSS nmos w=w_n l=lu

* Model comparator
*BC1 VCMP_OUT VSS V = ((atan(100000*(V(VSTORE) - V(VRAMP)))) + 1.58)/3.14*1.5


.ENDS
