* Current mirrors

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130.spi
.include ../../lib/SUN_TR_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-20


*----------------------------------------------------------------
* Paramater
.param w_n = 0.5u
.param w_p = {w_n * 2.57}
.param lu = 0.48u

* Sources 
VDD VDD VSS dc 1.5
VSS VSS 0 dc 0
V2 VSTORE 0 dc 0 
VRA VRAMP 0 dc 0.75
*----------------------------------------------------------------
* BIAS
*----------------------------------------------------------------
* Use a current mirror transistor from the SUN_TR_GF130N library
IPB1 0 VBN1 dc 1u
XMNB0 VBN1 VBN1 VSS VSS NCHCM2

* DUT
MP1 MPS1 MPS1 VDD VDD pmos w=w_p l=lu
MP2 MPS2 MPS1 VDD VDD pmos w=w_p l=lu
MN3 MPS1 VSTORE MNS3 MNS3 nmos w=w_n l=lu
MN4 MPS2 VRAMP MNS3 MNS3 nmos w=w_n l=lu
MN5 MNS3 VBN1 VSS VSS nmos w=w_n l=lu
MP6 MP6S MPS2 VDD VDD pmos w=w_p l=lu
MN7 MP6S VBN1 VSS VSS nmos w=w_n l=lu
MP8 TEST_OUT MP6S VDD VDD pmos w=w_p l=lu
MN9 TEST_OUT MP6S VSS VSS nmos w=w_n l=lu
MP10 VCMP_OUT TEST_OUT VDD VDD pmos w=w_p l=lu
MN11 VCMP_OUT TEST_OUT VSS VSS nmos w=w_n l=lu
* MN9 VCMP_OUT MP6S VSS VSS nmos w=w_n l=lu
*----------------------------------------------------------------
* Analysis
*----------------------------------------------------------------
.op
.dc V2 0.0 1.65 0.01
.plot dc V(V2) V(TEST_OUT) V(MNS3) V(VBN1)
 
